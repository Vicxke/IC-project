//------------------------------------------------------------------------------
//
// This module is a top-level module for the TB with serial data to parallel  DUT
//
// It instantiates all of the uVC interface instances and connects them to the RTL top.
// It also initializes the UVM test environment and runs the test and
// it creates the default top-level test configuration.
//
// The testbench uses the following uVC interfaces:
// - CLOCK IF: Generates a system clock.
// - RESET IF: Generates the reset signal.
// - SERIAL_DATA IF: Generate parallel data to the DUT input interface
// - PARALLEL_DATA IF: Passes the DUT output infterface to parallel data uVC
//
//------------------------------------------------------------------------------
module tb_top;

    // Include basic packages
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    import common::*;

    // Include optional packages
    import tb_pkg::*;

    // uVC TB signal variables
    logic tb_clock;
    logic tb_reset_n;

    // Instantiation of CLOCK uVC interface signal

    clock_if  i_clock_if();
    assign tb_clock = i_clock_if.clock;

    // Instantiation of RESET uVC interface signal
    reset_if  i_reset_if(.clk(tb_clock));
    assign tb_reset_n = i_reset_if.reset_n;

    // Instantiate execution_stage interface and connect to the DUT
    execution_stage_input_if i_execute_input_if(.clk(tb_clock), .rst_n(tb_reset_n));
    execution_stage_output_if i_execute_output_if(.clk(tb_clock), .rst_n(tb_reset_n));

    // decode stage interface instantiation would go here if needed
    decode_stage_input_if i_decode_input_if(.clk(tb_clock), .rst_n(tb_reset_n));

    decode_stage_output_if i_decode_output_if(.clk(tb_clock), .rst_n(tb_reset_n));


    // ------------------------------------------------------------
    // Declare signals that go from decode -> execute
    // (types must match your RTL ports!)
    // ------------------------------------------------------------
    logic [31:0] data1_decode_to_execute;
    logic [31:0] data2_decode_to_execute;
    logic [31:0] immediate_data_decode_to_execute;
    logic [31:0] program_counter_in_decode_to_execute;
    logic        compflg_in_decode_to_execute;
    control_type control_in_decode_to_execute; // from common::*
    bit          instr_valid_ex_in_decode_to_execute;

    
    // Instantiate decode_stage interface and connect to the DUT
    decode_stage dut_decode_stage (
        //inputs
        .clk(tb_clock),
        .reset_n(tb_reset_n),
        .instruction(i_decode_input_if.instruction),
        .pc(i_decode_input_if.pc),
        .compflg(i_decode_input_if.compflg),
        .write_en(i_decode_input_if.write_en),
        .write_id(i_decode_input_if.write_id),
        .write_data(i_decode_input_if.write_data),
        .mux_data1(i_decode_input_if.mux_data1),
        .mux_data2(i_decode_input_if.mux_data2),
        //outputs decode (no execution stage input)
        .reg_rd_id(i_decode_output_if.reg_rd_id),
        .select_target_pc(i_decode_output_if.select_target_pc),    //J-type is also taken into account
        .resolve(i_decode_output_if.resolve),                      //only high for B-type
        .squash_after_J(i_decode_output_if.squash_after_J), //sqaush from ID following a sequeatially fetched Jump
        .squash_after_JALR(i_decode_output_if.squash_after_JALR),
        .rs1_id(i_decode_output_if.rs1_id),
        .rs2_id(i_decode_output_if.rs2_id),

        // outputs decode inputs to execution stage
        .read_data1(data1_decode_to_execute),
        .read_data2(data2_decode_to_execute),
        .immediate_data(immediate_data_decode_to_execute),
        .control_signals(control_in_decode_to_execute),
        .calculated_target_pc(program_counter_in_decode_to_execute),
        .compflg_out(compflg_in_decode_to_execute)
    );

    
    // --------------------------------------------------------------------------
    // Wire DECODE outputs into the EXECUTE inputs (THIS is the critical part)
    // --------------------------------------------------------------------------
    assign i_execute_input_if.data1           = data1_decode_to_execute;
    assign i_execute_input_if.data2           = data2_decode_to_execute;
    assign i_execute_input_if.immediate_data  = immediate_data_decode_to_execute;
    assign i_execute_input_if.control_in      = control_in_decode_to_execute;
    assign i_execute_input_if.compflg_in      = compflg_in_decode_to_execute;
    assign i_execute_input_if.program_counter_in = program_counter_in_decode_to_execute;

    // pass instr_valid_ex_in from decode input interface to execute input and output interfaces
    assign i_execute_input_if.instr_valid_ex_in = i_decode_input_if.instr_valid_ex_in;
    assign i_execute_output_if.instr_valid_ex_in = i_decode_input_if.instr_valid_ex_in; 

    // pass instr_valid from decode input interface to decode output interface
    assign i_decode_output_if.instr_valid = i_decode_input_if.instr_valid;


    // Instantiation of the execute_stage RTL DUT
    execute_stage dut_execute_stage (
        //inputs
        .clk(tb_clock),
        .reset_n(tb_reset_n),
        .data1(i_execute_input_if.data1),
        .data2(i_execute_input_if.data2),
        .immediate_data(i_execute_input_if.immediate_data),
        .control_in(i_execute_input_if.control_in),
        .compflg_in(i_execute_input_if.compflg_in),
        .program_counter(i_execute_input_if.program_counter_in),
        //outpus
        .control_out(i_execute_output_if.control_out),
        .alu_data(i_execute_output_if.alu_data),
        .memory_data(i_execute_output_if.memory_data),
        .overflow_flag(i_execute_output_if.overflow_flag),
        .compflg_out(i_execute_output_if.compflg_out)
    );

    // --------------------- connection missing for decode stage DUT if applicable ---------------------
    always @(
        i_execute_input_if.data1,
        i_execute_input_if.data2,
        i_execute_input_if.immediate_data,
        i_execute_input_if.control_in,
        i_execute_input_if.program_counter_in,
        i_execute_input_if.compflg_in
    ) begin
        $display("[%0t] EX-IN:"
                , $time,
                " d1=%0h d2=%0h imm=%0h instr=%0h pc=%0h cmp=%0b",
                i_execute_input_if.data1,
                i_execute_input_if.data2,
                i_execute_input_if.immediate_data,
                i_execute_input_if.control_in.alu_op.name(),
                i_execute_input_if.program_counter_in,
                i_execute_input_if.compflg_in);       
    end


    always @(
        data1_decode_to_execute,
        data2_decode_to_execute,
        immediate_data_decode_to_execute,
        control_in_decode_to_execute,
        program_counter_in_decode_to_execute,
        compflg_in_decode_to_execute,
        i_decode_output_if.reg_rd_id
    ) begin
            $display("[%0t] DEC-OUT:"
                , $time,
                " d1=%0h d2=%0h imm=%0h instr=%0h pc=%0h cmp=%0b rd_id=%0h",
                data1_decode_to_execute,
                data2_decode_to_execute,
                immediate_data_decode_to_execute,
                control_in_decode_to_execute.alu_op.name(),
                program_counter_in_decode_to_execute,
                compflg_in_decode_to_execute,
                i_decode_output_if.reg_rd_id);       
    end

    always @(
        i_decode_input_if.instruction,
        i_decode_input_if.pc,
        i_decode_input_if.compflg,
        i_decode_input_if.write_en,
        i_decode_input_if.write_id,
        i_decode_input_if.write_data,
        i_decode_input_if.mux_data1,
        i_decode_input_if.mux_data2
    ) begin
            $display("[%0t] DEC-IN:"
                , $time,
                " instr=%0h pc=%0h comp=%0h write_en=%0h write_id=%0h write_data=%0h mux1=%0h mux2=%0h",
                i_decode_input_if.instruction,
                i_decode_input_if.pc,
                i_decode_input_if.compflg,
                i_decode_input_if.write_en,
                i_decode_input_if.write_id,
                i_decode_input_if.write_data,
                i_decode_input_if.mux_data1,
                i_decode_input_if.mux_data2);       
    end

    always @(
        i_execute_output_if.control_out,
        i_execute_output_if.alu_data,
        i_execute_output_if.memory_data,
        i_execute_output_if.overflow_flag,
        i_execute_output_if.compflg_out
    ) begin
            $display("[%0t] EXE-OUT:"
                , $time,
                " ctrl_out=%0h alu_data=%0h memory_data=%0h overflow_flag=%0h compflg_out=%0b",
                i_execute_output_if.control_out,
                i_execute_output_if.alu_data,
                i_execute_output_if.memory_data,
                i_execute_output_if.overflow_flag,
                i_execute_output_if.compflg_out);       
    end

    always @(
        i_execute_input_if.instr_valid_ex_in
    ) begin
        $display("[%0t] EX-INSTR_VALID:"
                , $time,
                " instr_valid_ex_in=%0b",
                i_execute_input_if.instr_valid_ex_in);       
    end


    // Initialize TB configuration
    initial begin
        top_config  m_top_config;
        // Create TB top configuration and store it into UVM config DB.
        m_top_config = new("m_top_config");
        uvm_config_db #(top_config)::set(null,"tb_top","top_config", m_top_config);
        // Save all virtual interface instances into configuration
        m_top_config.m_clock_config.m_vif = i_clock_if;
        m_top_config.m_reset_config.m_vif = i_reset_if;
        // Save execution_stage interface instance into top config
        m_top_config.m_execution_stage_input_config.m_vif = i_execute_input_if;
        m_top_config.m_execution_stage_output_config.m_vif = i_execute_output_if;
        // Save decode_stage interface instance into top config
        m_top_config.m_decode_stage_input_config.m_vif = i_decode_input_if;
        m_top_config.m_decode_stage_output_config.m_vif = i_decode_output_if;
    end

    // Start UVM test_base environment
    initial begin // only one run valid
        // run_test("ExDeStage_00"); 
        //run_test("ExDeStage_01"); 
        //run_test("ExDeStage_02"); 
        // run_test("ExDeStage_03");
        run_test("ExDeStage_04");
    end

endmodule
