//------------------------------------------------------------------------------
// Scoreboard for the TBUVM TB.
//
// This class is an implementation of the scoreboard that monitors the TBUVM
// testbench and checks the behavior of the DUT with regard to the
// serial-to-parallel conversion. It provides the following features:
//
// - Monitors the input serial data and the output parallel data of the DUT.
// - Checks if the output data of the DUT is correct with regard to the
//   input serial data.
// - Checks if the DUT is in the correct state during the transmission of data.
// - Provides functional coverage for the transmission of data and the
//   activation of the DUT's output.
// - Provides error reporting for any errors that are detected during the simulation.
//
// This class is derived from the `uvm_component` class and implements the
// `uvm_analysis_imp_scoreboard_reset`, `uvm_analysis_imp_scoreboard_serial_data`
// and `uvm_analysis_imp_scoreboard_parallel_data` analysis ports.
//
// The functional coverage is provided by the `serial_to_parallel_covergrp`
// coverage group.
//

import common::*;

//------------------------------------------------------------------------------
// Instance analysis defines (creates unique analysis_imp types)
`uvm_analysis_imp_decl(_scoreboard_reset)
`uvm_analysis_imp_decl(_scoreboard_execution_stage)

// Simplified scoreboard for execution_stage UVC
class scoreboard extends uvm_component;
    `uvm_component_utils(scoreboard)

    // execution_stage analysis connection (uses a dedicated analysis_imp type)
    uvm_analysis_imp_scoreboard_execution_stage#(execution_stage_seq_item, scoreboard) m_execution_stage_ap;
    // reset analysis connection
    uvm_analysis_imp_scoreboard_reset#(reset_seq_item, scoreboard) m_reset_ap;

    // basic counters
    int unsigned items_received = 0;

    // Indicates if the reset signal is active.
    //int unsigned reset_valid;
    // The value of the reset signal.
    int unsigned reset_value;
    // The ALU operation being performed.
    alu_op_type alu_op;

    int unsigned data1;
    int unsigned data2;

    encoding_type encoding;

    //------------------------------------------------------------------------------
    // Functional coverage definitions
    //------------------------------------------------------------------------------
    covergroup execution_stage_covergrp;
        reset : coverpoint reset_value {
            bins reset =  { 0 };
            bins run=  { 1 };
        }
        operations : coverpoint alu_op {
            bins ADD =  { ALU_ADD };
            bins SUB =  { ALU_SUB };
            bins XOR =  { ALU_XOR };
            bins OR  =  { ALU_OR };
            bins AND =  { ALU_AND };
            bins SLL =  { ALU_SLL };
            bins SRL =  { ALU_SRL };
            bins SRA =  { ALU_SRA };
            bins SLT =  { ALU_SLT };
            bins SLTU=  { ALU_SLTU };
        }
        operand_1 : coverpoint data1 {
            bins very_low   = { [32'h00000000 : 32'h0000FFFF] };   
            bins low        = { [32'h00010000 : 32'h00FFFFFF] };    
            bins mid_low    = { [32'h01000000 : 32'h0FFFFFFF] };    
            bins mid        = { [32'h10000000 : 32'h3FFFFFFF] };   
            bins mid_high   = { [32'h40000000 : 32'h7FFFFFFF] };   
            bins high       = { [32'h80000000 : 32'hBFFFFFFF] };   
            bins very_high  = { [32'hC0000000 : 32'hEFFFFFFF] };    
            bins max_val    = { [32'hF0000000 : 32'hFFFFFFFF] };     
        }
        operand_2 : coverpoint data2 {
            bins very_low   = { [32'h00000000 : 32'h0000FFFF] };   
            bins low        = { [32'h00010000 : 32'h00FFFFFF] };    
            bins mid_low    = { [32'h01000000 : 32'h0FFFFFFF] };    
            bins mid        = { [32'h10000000 : 32'h3FFFFFFF] };   
            bins mid_high   = { [32'h40000000 : 32'h7FFFFFFF] };   
            bins high       = { [32'h80000000 : 32'hBFFFFFFF] };   
            bins very_high  = { [32'hC0000000 : 32'hEFFFFFFF] };    
            bins max_val    = { [32'hF0000000 : 32'hFFFFFFFF] };     
        }
        op_type : coverpoint encoding {
            bins R_TYPE = { R_TYPE };
            bins I_TYPE = { I_TYPE };
            bins S_TYPE = { S_TYPE };
            bins B_TYPE = { B_TYPE };
            bins U_TYPE = { U_TYPE };
            bins J_TYPE = { J_TYPE };
        }
        cross_op_reset : cross operations, reset; //test cross coverage
        cross_op_data : cross operations, operand_1, operand_2;
    endgroup

    //------------------------------------------------------------------------------
    // The constructor for the component.
    //------------------------------------------------------------------------------
    function new(string name = "scoreboard", uvm_component parent = null);
        super.new(name,parent);
        // Create coverage group
        execution_stage_covergrp = new();
    endfunction: new

    //------------------------------------------------------------------------------
    // The build for the component.
    //------------------------------------------------------------------------------
    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        m_execution_stage_ap = new("m_execution_stage_ap", this);
        m_reset_ap = new("m_reset_ap", this);
    endfunction: build_phase

    //------------------------------------------------------------------------------
    // The connection phase for the component.
    //------------------------------------------------------------------------------
    virtual function void connect_phase(uvm_phase phase);
        super.connect_phase(phase);
    endfunction: connect_phase

    //------------------------------------------------------------------------------
    // Write implementation for write_scoreboard_execution_stage analysis port.
    //------------------------------------------------------------------------------
    virtual function void write_scoreboard_execution_stage(execution_stage_seq_item item);
        `uvm_info(get_name(), $sformatf("EXECUTION_STAGE_MONITOR: %s", item.convert2string()), UVM_MEDIUM)
        items_received++;
        if (item.exp_alu_data !== 'x && item.exp_alu_data !== '0) begin
            `uvm_info(get_name(), $sformatf("Item provided expected ALU data=0x%08h", item.exp_alu_data), UVM_LOW)
        end

        alu_op= item.control_in.alu_op;
        data1 = item.data1;
        data2 = item.data2;
        encoding = item.control_in.encoding;
        //`uvm_info(get_name(), $sformatf("ALU_OPRESET_function: alu_op=%00s reset_value=%0b", alu_op.name(), reset_value), UVM_LOW)
        execution_stage_covergrp.sample();

    endfunction: write_scoreboard_execution_stage

    //------------------------------------------------------------------------------
    // Write implementation for write_scoreboard_reset analysis port.
    //------------------------------------------------------------------------------
    virtual function void write_scoreboard_reset(reset_seq_item item);
        `uvm_info(get_name(),$sformatf("RESET_MONITOR:\n%s",item.sprint()),UVM_HIGH)
        // // Clear start bit and data
        // input_data_valid= 0;
        // input_data= 0;
        // dut_data_valid= 0;
        // dut_data= 0;
        // Sample reset coverage
        reset_value= item.reset_value;
        //`uvm_info(get_name(), $sformatf("RESET_function: alu_op=%00s reset_value=%0b", alu_op.name(), reset_value), UVM_LOW)
        execution_stage_covergrp.sample();

    endfunction :  write_scoreboard_reset

    //------------------------------------------------------------------------------
    // UVM check phase
    //------------------------------------------------------------------------------
    virtual function void check_phase(uvm_phase phase);
        super.check_phase(phase);
        $display("*****************************************************");
        if (execution_stage_covergrp.get_coverage() == 100.0) begin
            $display("FUNCTIONAL COVERAGE (100.0%%) PASSED....");
        end
        else begin
            $display("FUNCTIONAL COVERAGE FAILED!!!!!!!!!!!!!!!!!");
            $display("Coverage = %0f", execution_stage_covergrp.get_coverage());
        end
        $display("*****************************************************");
    endfunction : check_phase

endclass: scoreboard
